ENTITY calculadora IS 
	PORT(
		XE1,XE2:IN BIT_VECTOR(3 DOWNTO 0);
		Sm2,Sm1,Sm0,BLigar:IN BIT;
		SaidaDisplay:OUT BIT_VECTOR(6 DOWNTO 0);
		LED:OUT BIT);
END calculadora;
ARCHITECTURE converteDisplay OF calculadora IS
COMPONENT SOMA4BITS 
	PORT(Carryin:IN BIT;
		X1,X2:IN BIT_VECTOR(3 DOWNTO 0);
		Sout:OUT BIT_VECTOR(3 DOWNTO 0);
	Carryout:OUT BIT);
END COMPONENT;
COMPONENT DECODIFICADORDISPLAY 
	PORT(
		CONTRL:IN BIT;
		ED:IN BIT_VECTOR(3 DOWNTO 0);
		VetorSaida:OUT BIT_VECTOR(6 DOWNTO 0));
END COMPONENT;
COMPONENT MULTIPLEXADOR4BITS
		PORT(
		Em14B,Em24B,Em34B,Em44B:IN BIT_VECTOR(3 DOWNTO 0);
		Em11B,Em21B,Em31B,Em41B,Em51B,Em61B:IN BIT;
		S01,S11,S21,BLD:IN BIT;
		VetorSaida:OUT BIT_VECTOR(3 DOWNTO 0);
		Cout,Ctrl:OUT BIT);
END COMPONENT;
COMPONENT COMPARADOR4BITS 
	PORT(
		SE41,SE42:BIT_VECTOR(3 DOWNTO 0);
		SE4q,SM4t,SL4t:OUT BIT);
END COMPONENT;
COMPONENT SUBTRACAOC2  
	PORT(
		SE1,SE2:IN BIT_VECTOR(3 DOWNTO 0);
		SUBOut:OUT BIT_VECTOR(3 DOWNTO 0);
		SignOut:OUT BIT);
END COMPONENT;
COMPONENT INVERSORC2 
	PORT(
		EC21:IN BIT_VECTOR(3 DOWNTO 0);
		nC2E:OUT BIT_VECTOR(3 DOWNTO 0);
	Cout:OUT BIT);
END COMPONENT;
COMPONENT INVERSORB  
	PORT(
		E1:IN BIT_VECTOR(3 DOWNTO 0);
		nE:OUT BIT_VECTOR(3 DOWNTO 0));
END COMPONENT;
SIGNAL Som:BIT_VECTOR(3 DOWNTO 0);
SIGNAL Sub:BIT_VECTOR(3 DOWNTO 0);
SIGNAL INVC2:BIT_VECTOR(3 DOWNTO 0);
SIGNAL INV:BIT_VECTOR(3 DOWNTO 0);
SIGNAL SAIDAMUX:BIT_VECTOR(3 DOWNTO 0); 
SIGNAL CARRY:BIT_VECTOR(5 DOWNTO 0);
SIGNAL Control:BIT;
BEGIN
SOMA: SOMA4BITS PORT MAP(Carryin=>'0',X1=>XE1,X2=>XE2,Sout=>Som,Carryout=>CARRY(0));
SUBTRACAO:SUBTRACAOC2 PORT MAP(SE1=>XE1,SE2=>XE2,SUBOut=>Sub,SignOut=>CARRY(1));
INVERSO: INVERSORB PORT MAP(E1=>XE1,nE=>INV);
INVERSOC2: INVERSORC2 PORT MAP(EC21=>XE1,nC2E=>INVC2,Cout=>CARRY(2));
COMPARACAO:COMPARADOR4BITS PORT MAP(SE41=>XE1,SE42=>XE2,SE4q=>CARRY(3),SM4t=>CARRY(4),SL4t=>CARRY(5));
MUX: MULTIPLEXADOR4BITS PORT MAP(Em14B=>Som,Em24B=>Sub,Em34B=>INV,Em44B=>INVC2,Em11B=>CARRY(0),Em21B=>CARRY(1),Em31B=>'0',Em41B=>CARRY(2),Em51B=>CARRY(4),Em61B=>CARRY(5),S01=>Sm0,S11=>Sm1,S21=>Sm2,BLD=>BLigar,VetorSaida=>SAIDAMUX,Cout=>LED,Ctrl=>Control);
DISPLAY7SEG: DECODIFICADORDISPLAY PORT MAP(CONTRL=>Control,ED=>SAIDAMUX,VetorSaida=>SAIdaDisplay);
END converteDisplay;
