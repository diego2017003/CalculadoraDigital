ENTITY COMPARADOR4BITS IS 
	PORT(
		SE41,SE42:BIT_VECTOR(3 DOWNTO 0);
		SE4q,SM4t,SL4t:OUT BIT);
END COMPARADOR4BITS;
ARCHITECTURE compara4BIT OF COMPARADOR4BITS IS
COMPONENT COMPARADOR1BIT 
PORT(
		SE1,SE2,SoEq,SoMt,SoLt:IN BIT;
		SEq,SMt,SLt:OUT BIT);
END COMPONENT;
SIGNAL S1:BIT_VECTOR(11 DOWNTO 0);
BEGIN
	C:COMPARADOR1BIT PORT MAP(SE1=>SE41(3),SE2=>SE42(3),SoEq=>'1',SoMt=>'0',SoLt=>'0',SEq=>S1(0),SMt=>S1(1),SLt=>S1(2));
	C2:COMPARADOR1BIT PORT MAP(SE1=>SE41(2),SE2=>SE42(2),SoEq=>S1(0),SoMt=>S1(1),SoLt=>S1(2),SEq=>S1(3),SMt=>S1(4),SLt=>S1(5));
	C3:COMPARADOR1BIT PORT MAP(SE1=>SE41(1),SE2=>SE42(1),SoEq=>S1(3),SoMt=>S1(4),SoLt=>S1(5),SEq=>S1(6),SMt=>S1(7),SLt=>S1(8));
	C4:COMPARADOR1BIT PORT MAP(SE1=>SE41(0),SE2=>SE42(0),SoEq=>S1(6),SoMt=>S1(7),SoLt=>S1(8),SEq=>S1(9),SMt=>S1(10),SLt=>S1(11));

	SE4q<=S1(9);
	SM4t<=S1(10);
	SL4t<=S1(11);
END compara4BIT;
