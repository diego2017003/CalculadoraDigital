ENTITY SUBTRACAOC2 IS 
	PORT(
		SE1,SE2:IN BIT_VECTOR(3 DOWNTO 0);
		SUBOut:OUT BIT_VECTOR(3 DOWNTO 0);
		SignOut:OUT BIT);
END SUBTRACAOC2;
ARCHITECTURE subtraic2 OF SUBTRACAOC2 IS
COMPONENT SOMA4BITS
	PORT(Carryin:IN BIT;
		X1,X2:IN BIT_VECTOR(3 DOWNTO 0);
		Sout:OUT BIT_VECTOR(3 DOWNTO 0);
	Carryout:OUT BIT);
END COMPONENT;
COMPONENT INVERSORB
	PORT(
		E1:IN BIT_VECTOR(3 DOWNTO 0);
		nE:OUT BIT_VECTOR(3 DOWNTO 0));
END COMPONENT;
SIGNAL INV:BIT_VECTOR(3 DOWNTO 0);
BEGIN
	INVERTEE2:INVERSORB PORT MAP(E1=>SE2,nE=>INV);
	subtracao:SOMA4BITS PORT MAP(Carryin=>'1',X1=>SE1,X2=>INV,Sout=>SUBOut,Carryout=>SignOut);
END subtraic2;
