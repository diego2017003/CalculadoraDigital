ENTITY INVERSORB IS 
	PORT(
		E1:IN BIT_VECTOR(3 DOWNTO 0);
		nE:OUT BIT_VECTOR(3 DOWNTO 0));
END INVERSORB;
ARCHITECTURE inverte OF INVERSORB IS
BEGIN
	nE(0)<=NOT(E1(0));
	nE(1)<=NOT(E1(1));
	nE(2)<=NOT(E1(2));
	nE(3)<=NOT(E1(3));
END inverte;
