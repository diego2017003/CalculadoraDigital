ENTITY DECODIFICADORDISPLAY IS 
	PORT(
		CONTRL:IN BIT;
		ED:IN BIT_VECTOR(3 DOWNTO 0);
		VetorSaida:OUT BIT_VECTOR(6 DOWNTO 0));
END DECODIFICADORDISPLAY;
ARCHITECTURE converteDisplay OF DECODIFICADORDISPLAY IS
SIGNAL INTERM:BIT_VECTOR(6 DOWNTO 0);
BEGIN
INTERM(0)<=((ED(3) XNOR ED(2))AND(NOT(ED(1)))AND((ED(0))))OR((NOT(ED(3)))AND(ED(2))AND(NOT(ED(1)))AND(NOT(ED(0))))OR((ED(3))AND(NOT(ED(2))AND(ED(1))AND(ED(0)))); 
INTERM(1)<=(ED(1)AND(ED(2))AND(NOT(ED(0))))OR(ED(3)AND(ED(2))AND(NOT(ED(0))))OR(ED(1)AND(ED(3))AND(ED(0)))OR((NOT ED(1))AND(ED(2))AND(ED(0))AND(NOT(ED(3))));
INTERM(2)<=((NOT ED(3))AND(ED(1))AND(NOT ED(2))AND(NOT(ED(0))))OR((ED(3))AND(ED(2))AND((ED(1))OR(NOT ED(0))));
INTERM(3)<=(ED(0)AND((ED(1)AND(ED(2)))OR((NOT ED(1))AND(NOT ED(2))AND(NOT(ED(3))))))OR((NOT ED(0))AND(((ED(1))AND((NOT ED(2))AND((ED(3)))))OR((NOT ED(1))AND(ED(2))AND(NOT(ED(3))))));
INTERM(4)<=(ED(0)AND((NOT(ED(3)))OR((NOT ED(2))AND(NOT ED(1)))))OR((NOT ED(3))AND(ED(2))AND(NOT ED(1)));
INTERM(5)<=((NOT ED(3))AND(NOT ED(2))AND(ED(1) OR ED(0)))OR(ED(0)AND(((NOT ED(3))AND(ED(1)))OR((ED(3))AND(ED(2))AND(NOT ED(1)))));
INTERM(6)<=((NOT ED(3))AND(((NOT ED(2))AND(NOT ED(1)))OR((ED(2))AND(ED(1))AND(ED(0)))))OR((ED(3))AND(ED(2))AND(NOT ED(1))AND(NOT ED(0)));

vetorSaida(0)<=(CONTRL AND INTERM(0))OR(NOT CONTRL);
vetorSaida(1)<=(CONTRL AND INTERM(1))OR(NOT CONTRL);
vetorSaida(2)<=(CONTRL AND INTERM(2))OR(NOT CONTRL);
vetorSaida(3)<=(CONTRL AND INTERM(3))OR(NOT CONTRL);
vetorSaida(4)<=(CONTRL AND INTERM(4))OR(NOT CONTRL);
vetorSaida(5)<=(CONTRL AND INTERM(5))OR(NOT CONTRL);
vetorSaida(6)<=(CONTRL AND INTERM(6))OR(NOT CONTRL);

END converteDisplay;
